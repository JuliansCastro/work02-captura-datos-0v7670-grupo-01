`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:27:31 11/12/2019 
// Design Name: 
// Module Name:    Captura 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Captura(
    input [7:0] Data,
    input Href,
    input Vsync,
    input Pclk,
    output regWrite,
    output addr_in
    );


endmodule
